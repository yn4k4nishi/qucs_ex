module logicgate_or( A, Y, B ) ;
	input A, B ;
	output Y ;
	assign Y = A | B ;
endmodule